version https://git-lfs.github.com/spec/v1
oid sha256:31fa019f2d8840213b3e64fb4468fb67e810f2016f7e4da46b005814675d7a37
size 80831540
