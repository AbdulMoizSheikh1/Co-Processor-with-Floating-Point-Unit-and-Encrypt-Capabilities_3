version https://git-lfs.github.com/spec/v1
oid sha256:135ba7d1e5e6b615dfaaf8466009e7e41f040579cdcb0a803db1f5b5cee95c00
size 169377
