version https://git-lfs.github.com/spec/v1
oid sha256:2f65c3bfad4e4c34ab2f325063d0e383bb0e76a44d902f5d09740e6330699eac
size 131256
