version https://git-lfs.github.com/spec/v1
oid sha256:1c0ba96eb30658128cf8e14af49157a6023e6dddea5a3b3a290c7a214da2bedc
size 3433539
